`include "defines.v"

module ROB(

    //output
    output wire             enCDBWrt, 
    output wire[`NameBus]   CDBwrtName, 
    output wire[`TagBus]    CDBwrtTag, 
    output wire[`DataBus]   CDBwrtData
)

endmodule
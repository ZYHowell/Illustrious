`include "defines.v"

module fetch(

)

endmodule